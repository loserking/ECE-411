import lc3b_types::*;

module mp3
(
    input clk

);

/* Instantiate MP 3 top level blocks here */



endmodule : mp3
