/*calculates and*/

module and2input(
		input logic x, y,
		output logic z
		
);

assign z = x & y;

endmodule : and2input