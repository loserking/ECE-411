/*calculates and*/

module or2input(
		input wire x, y,
		output wire z
		
);

assign z = x | y;

endmodule : or2input