/*calculates and*/

module and2input(
		input wire x, y,
		output wire z
		
);

assign z = x & y;

endmodule : and2input